module topl(
    parameter ADDRESS_WIDTH=5,
              DATA_WIDTH=32
)(

    input logic clk,
    input logic RegWrite,
    input 
)
;


endmodule