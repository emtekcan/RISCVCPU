module simplecpu(
    input logic clk,
    input logic rst
);

pcreg PC(


);

cutop CU(


);

alutop ALU(


);





endmodule